//========================================================================== //
// Copyright (c) 2026, Stephen Henry
// All rights reserved.
//
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// * Redistributions of source code must retain the above copyright notice, this
//   list of conditions and the following disclaimer.
//
// * Redistributions in binary form must reproduce the above copyright notice,
//   this list of conditions and the following disclaimer in the documentation
//   and/or other materials provided with the distribution.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
// ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
// INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
// CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.
//========================================================================== //

`include "common_defs.svh"
`include "math_pkg.svh"

// Circuit to compute the cicular left-most '0' in a vector 'x' for a
// given position. 'any' flag indicates output validity.
//
//   x                       pos   y                      y_enc    any
//   -----------------------------------------------------------------------
//
//   1111_1111_1111_1110     0     0000_0000_0000_0001    0        1
//                     ^
//
//   0000_0000_0000_0000     0     1000_0000_0000_0000    15       1
//                     ^
//
//   0000_0000_0000_0000     1     0000_0000_0000_0001    0        1
//                    ^
//
//   0000_0000_0000_0000    15     0100_0000_0000_0000    14       1
//   ^
//
//   0010_1010_0011_0111     8     0000_0000_1000_0000    7        1
//           ^
//
//   1111_1111_1111_1111     x     xxxx_xxxx_xxxx_xxxx    x        0

module e_multi #(
  // Vector width
  parameter int W = 32

  // Radix (In range: [4,8])
, parameter int RADIX_N = 4
) (
  input wire logic [W - 1:0]                     x_i
, input wire logic [$clog2(W) - 1:0]             pos_i

//
, output wire logic [W - 1:0]                    y_o
, output wire logic [$clog2(W) - 1:0]            y_enc_o
, output wire logic                              any_o
);

// ========================================================================= //
//                                                                           //
// Localparams                                                               //
//                                                                           //
// ========================================================================= //

localparam int SEARCH_WORD_W = 2 * W;

localparam int GROUPS_N = math_pkg::div_ceil(SEARCH_WORD_W, RADIX_N);

typedef logic [GROUPS_N - 1:0]                     groups_t;
typedef logic [GROUPS_N - 1:0][RADIX_N - 1:0]      groups_vec_t;

localparam int GROUPS_VEC_W = $bits(groups_vec_t);

// Flag indicating whether the groups require padding to fill the last group.
localparam bit REQUIRES_PADDING = (GROUPS_N * RADIX_N != SEARCH_WORD_W);


// ========================================================================= //
//                                                                           //
// Wire(s)                                                                   //
//                                                                           //
// ========================================================================= //

logic [W - 1:0]                        pos_dec;

groups_t                               groups_prior;
groups_vec_t                           groups_sel;
groups_vec_t                           groups_in;
groups_vec_t                           groups_out;
groups_t                               groups_out_vld;

logic                                  any;

logic [W - 1:0]                        y;
logic [$clog2(W) - 1:0]                y_enc;

// ========================================================================= //
//                                                                           //
// Logic.                                                                    //
//                                                                           //
// ========================================================================= //

// ------------------------------------------------------------------------- //
// Compute selection vector.
dec #(.W(W)) u_dec (
  .x_i                       (pos_i)
, .y_o                       (pos_dec)
);

// ------------------------------------------------------------------------- //
// Compute input vector (padding if required).
if (REQUIRES_PADDING) begin : gen_groups_padding
  localparam int PADDING_BITS = (GROUPS_N * RADIX_N) - W;

  assign groups_in = { {(PADDING_BITS{1'b0}}, x_i, x_i };
  assign groups_sel = { {(PADDING_BITS{1'b0}}, pos_dec, pos_dec };
end
else begin : gen_groups_no_padding

  assign groups_in = { x_i, x_i };
  assign groups_sel = { pos_dec, pos_dec };
end : gen_groups_no_padding

// ------------------------------------------------------------------------- //
// Groups prior:
for (genvar i = 0; i < GROUPS_N; i++) begin : group_prior_GEN

if (i == (GROUPS_N - 1)) begin: last_group_GEN

  assign groups_prior[i] = 1'b0;
end: last_group_GEN
else begin: not_last_group_GEN
  localparam int j = (i * RADIX_N);

  assign groups_prior[i] = (groups_in[j] & groups_sel[j]);
end: not_last_group_GEN

end : group_prior_GEN

// ------------------------------------------------------------------------- //
//
for (genvar i = 0; i < GROUPS_N; i++) begin : group_GEN

  e_priority #(.W(RADIX_N)) u_e_priority (
    .x_prior_and_sel_i       (groups_prior[i])
  , .x_i                     (groups_in[i])
  , .sel_i                   (groups_sel[i])
  , .vld_o                   (groups_out_vld[i])
  , .y_o                     (groups_out[i]));

end : group_GEN

// ------------------------------------------------------------------------- //
//
for (genvar i = 0; i < GROUPS_N; i++) begin: group_cell_GEN

if (i == (GROUPS_N - 1)) begin: last_group_cell_GEN

  e_multi_cell u_e_multi_cell (
    .vld_i                    (groups_out_vld[i])
  , .prior_i                  (1'b0)
  , .sel_i                    (groups_sel[(i * RADIX_N) +: RADIX_N])
  //
  , .next_o                   ()
  );

  end: last_group_cell_GEN

else begin: not_last_group_cell_GEN

  e_multi_cell u_e_multi_cell (
    .vld_i                    (groups_out_vld[i])
  , .prior_i                  (1'b0)
  , .sel_i                    (groups_sel[(i * RADIX_N) +: RADIX_N])
  //
  , .next_o                   ()
  );

end: group_cell_GEN

// ------------------------------------------------------------------------- //
// If no bit is found in the bits preceeding pos_i, use the output
// from the succeeding bits logic.
//
assign y = '0;


// ------------------------------------------------------------------------- //
// 'Any' flag; indicate that a 'b0 is present in the input vector. The
// output at y_* is therefore valid.
// 
assign any = (x_i != '1);


// ------------------------------------------------------------------------- //
// Compute encoded output.
enc #(.W(W)) u_enc (.x_i(y), .y_o(y_enc));


// ========================================================================= //
//                                                                           //
// Output(s)                                                                 //
//                                                                           //
// ========================================================================= //

assign any_o = any;
assign y_o = y;
assign y_enc_o = y_enc;

endmodule : e_multi
